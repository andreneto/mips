module cpu();
endmodule