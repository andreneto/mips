module cpu(clock);
endmodule