module mult(in_0, in_1, out_0, out_1);
input wire [31:0] in_0, in_1;
output reg [31:0] out_0, out_1;


endmodule